

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity xor_gate2 is
	port(A : in std_logic;
			B : in std_logic;
			Y : out std_logic;
			);
end xor_gate2




