module xor_gate_test (
    input A,
    input B,
    output Y
);
    assign Y = A ^ B;
endmodule
